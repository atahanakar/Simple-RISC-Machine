module shifter #(
    data_width = 16
  )(
    // INPUTS
    input logic  [data_width - 1:0] in,
    input logic  [1:0] shift,
    // OUTPUTS
    output logic [data_width - 1:0] sout1
  );
  // Insert the code here

endmodule
