module ALU(
  parameter data_width = 16
  )(
  // INPUTS
  input logic  [data_width - 1:0] Ain,
  input logic  [data_width - 1:0] Bin,

  // OUTPUTS
  output logic [data_width - 1:0] out,
  output logic Z
  );


endmodule
